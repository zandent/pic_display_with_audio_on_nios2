
module sub_top (
	clk_clk,
	reset_reset_n,
	audio_0_external_interface_BCLK,
	audio_0_external_interface_DACDAT,
	audio_0_external_interface_DACLRCK);	

	input		clk_clk;
	input		reset_reset_n;
	input		audio_0_external_interface_BCLK;
	output		audio_0_external_interface_DACDAT;
	input		audio_0_external_interface_DACLRCK;
endmodule
