// sub_top.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module sub_top (
		input  wire        audio_0_external_interface_BCLK,                 //                audio_0_external_interface.BCLK
		output wire        audio_0_external_interface_DACDAT,               //                                          .DACDAT
		input  wire        audio_0_external_interface_DACLRCK,              //                                          .DACLRCK
		input  wire        clk_clk,                                         //                                       clk.clk
		output wire [12:0] new_sdram_controller_0_wire_addr,                //               new_sdram_controller_0_wire.addr
		output wire [1:0]  new_sdram_controller_0_wire_ba,                  //                                          .ba
		output wire        new_sdram_controller_0_wire_cas_n,               //                                          .cas_n
		output wire        new_sdram_controller_0_wire_cke,                 //                                          .cke
		output wire        new_sdram_controller_0_wire_cs_n,                //                                          .cs_n
		inout  wire [15:0] new_sdram_controller_0_wire_dq,                  //                                          .dq
		output wire [1:0]  new_sdram_controller_0_wire_dqm,                 //                                          .dqm
		output wire        new_sdram_controller_0_wire_ras_n,               //                                          .ras_n
		output wire        new_sdram_controller_0_wire_we_n,                //                                          .we_n
		input  wire        reset_reset_n,                                   //                                     reset.reset_n
		output wire        video_vga_controller_0_external_interface_CLK,   // video_vga_controller_0_external_interface.CLK
		output wire        video_vga_controller_0_external_interface_HS,    //                                          .HS
		output wire        video_vga_controller_0_external_interface_VS,    //                                          .VS
		output wire        video_vga_controller_0_external_interface_BLANK, //                                          .BLANK
		output wire        video_vga_controller_0_external_interface_SYNC,  //                                          .SYNC
		output wire [7:0]  video_vga_controller_0_external_interface_R,     //                                          .R
		output wire [7:0]  video_vga_controller_0_external_interface_G,     //                                          .G
		output wire [7:0]  video_vga_controller_0_external_interface_B      //                                          .B
	);

	wire         video_dma_controller_0_avalon_pixel_source_valid;                             // video_dma_controller_0:stream_valid -> video_vga_controller_0:valid
	wire  [29:0] video_dma_controller_0_avalon_pixel_source_data;                              // video_dma_controller_0:stream_data -> video_vga_controller_0:data
	wire         video_dma_controller_0_avalon_pixel_source_ready;                             // video_vga_controller_0:ready -> video_dma_controller_0:stream_ready
	wire         video_dma_controller_0_avalon_pixel_source_startofpacket;                     // video_dma_controller_0:stream_startofpacket -> video_vga_controller_0:startofpacket
	wire         video_dma_controller_0_avalon_pixel_source_endofpacket;                       // video_dma_controller_0:stream_endofpacket -> video_vga_controller_0:endofpacket
	wire         sys_sdram_pll_0_sdram_clk_clk;                                                // sys_sdram_pll_0:sdram_clk_clk -> [audio_0:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_1:sys_sdram_pll_0_sdram_clk_clk, new_sdram_controller_0:clk, nios2_qsys_0:clk, onchip_memory2_0:clk, rst_controller:clk]
	wire         sys_sdram_pll_0_sys_clk_clk;                                                  // sys_sdram_pll_0:sys_clk_clk -> [avalon_MM_4_to_1_adapter_0:clock, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, mm_interconnect_1:sys_sdram_pll_0_sys_clk_clk, rst_controller_001:clk, video_dma_controller_0:clk, video_vga_controller_0:clk]
	wire         sys_sdram_pll_0_reset_source_reset;                                           // sys_sdram_pll_0:reset_source_reset -> [avalon_MM_4_to_1_adapter_0:reset_n, rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire         video_dma_controller_0_avalon_dma_master_waitrequest;                         // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_waitrequest -> video_dma_controller_0:master_waitrequest
	wire  [31:0] video_dma_controller_0_avalon_dma_master_readdata;                            // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdata -> video_dma_controller_0:master_readdata
	wire  [31:0] video_dma_controller_0_avalon_dma_master_address;                             // video_dma_controller_0:master_address -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_address
	wire         video_dma_controller_0_avalon_dma_master_read;                                // video_dma_controller_0:master_read -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_read
	wire         video_dma_controller_0_avalon_dma_master_readdatavalid;                       // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdatavalid -> video_dma_controller_0:master_readdatavalid
	wire         video_dma_controller_0_avalon_dma_master_lock;                                // video_dma_controller_0:master_arbiterlock -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_lock
	wire  [31:0] mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_readdata;           // avalon_MM_4_to_1_adapter_0:s_readdata -> mm_interconnect_0:avalon_MM_4_to_1_adapter_0_avalon_slave_readdata
	wire         mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_waitrequest;        // avalon_MM_4_to_1_adapter_0:s_waitrequest -> mm_interconnect_0:avalon_MM_4_to_1_adapter_0_avalon_slave_waitrequest
	wire  [26:0] mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_address;            // mm_interconnect_0:avalon_MM_4_to_1_adapter_0_avalon_slave_address -> avalon_MM_4_to_1_adapter_0:s_address
	wire         mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_read;               // mm_interconnect_0:avalon_MM_4_to_1_adapter_0_avalon_slave_read -> avalon_MM_4_to_1_adapter_0:s_read
	wire         mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_readdatavalid;      // avalon_MM_4_to_1_adapter_0:s_readdatavalid -> mm_interconnect_0:avalon_MM_4_to_1_adapter_0_avalon_slave_readdatavalid
	wire         mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_lock;               // mm_interconnect_0:avalon_MM_4_to_1_adapter_0_avalon_slave_lock -> avalon_MM_4_to_1_adapter_0:s_lock
	wire         avalon_mm_4_to_1_adapter_0_avalon_master_chipselect;                          // avalon_MM_4_to_1_adapter_0:m_chipselect -> mm_interconnect_1:avalon_MM_4_to_1_adapter_0_avalon_master_chipselect
	wire         avalon_mm_4_to_1_adapter_0_avalon_master_waitrequest;                         // mm_interconnect_1:avalon_MM_4_to_1_adapter_0_avalon_master_waitrequest -> avalon_MM_4_to_1_adapter_0:m_waitrequest
	wire  [15:0] avalon_mm_4_to_1_adapter_0_avalon_master_readdata;                            // mm_interconnect_1:avalon_MM_4_to_1_adapter_0_avalon_master_readdata -> avalon_MM_4_to_1_adapter_0:m_readdata
	wire  [26:0] avalon_mm_4_to_1_adapter_0_avalon_master_address;                             // avalon_MM_4_to_1_adapter_0:m_address -> mm_interconnect_1:avalon_MM_4_to_1_adapter_0_avalon_master_address
	wire   [1:0] avalon_mm_4_to_1_adapter_0_avalon_master_byteenable;                          // avalon_MM_4_to_1_adapter_0:m_byteenable -> mm_interconnect_1:avalon_MM_4_to_1_adapter_0_avalon_master_byteenable
	wire         avalon_mm_4_to_1_adapter_0_avalon_master_read;                                // avalon_MM_4_to_1_adapter_0:m_read -> mm_interconnect_1:avalon_MM_4_to_1_adapter_0_avalon_master_read
	wire         avalon_mm_4_to_1_adapter_0_avalon_master_readdatavalid;                       // mm_interconnect_1:avalon_MM_4_to_1_adapter_0_avalon_master_readdatavalid -> avalon_MM_4_to_1_adapter_0:m_readdatavalid
	wire         avalon_mm_4_to_1_adapter_0_avalon_master_lock;                                // avalon_MM_4_to_1_adapter_0:m_lock -> mm_interconnect_1:avalon_MM_4_to_1_adapter_0_avalon_master_lock
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                            // mm_interconnect_1:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                                         // mm_interconnect_1:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                                         // nios2_qsys_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_qsys_0_data_master_debugaccess
	wire  [26:0] nios2_qsys_0_data_master_address;                                             // nios2_qsys_0:d_address -> mm_interconnect_1:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                          // nios2_qsys_0:d_byteenable -> mm_interconnect_1:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                                // nios2_qsys_0:d_read -> mm_interconnect_1:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                                               // nios2_qsys_0:d_write -> mm_interconnect_1:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                           // nios2_qsys_0:d_writedata -> mm_interconnect_1:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                                     // mm_interconnect_1:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                                  // mm_interconnect_1:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [13:0] nios2_qsys_0_instruction_master_address;                                      // nios2_qsys_0:i_address -> mm_interconnect_1:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                                         // nios2_qsys_0:i_read -> mm_interconnect_1:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_1_new_sdram_controller_0_s1_chipselect;                       // mm_interconnect_1:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire  [15:0] mm_interconnect_1_new_sdram_controller_0_s1_readdata;                         // new_sdram_controller_0:za_data -> mm_interconnect_1:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_1_new_sdram_controller_0_s1_waitrequest;                      // new_sdram_controller_0:za_waitrequest -> mm_interconnect_1:new_sdram_controller_0_s1_waitrequest
	wire  [24:0] mm_interconnect_1_new_sdram_controller_0_s1_address;                          // mm_interconnect_1:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_1_new_sdram_controller_0_s1_read;                             // mm_interconnect_1:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire   [1:0] mm_interconnect_1_new_sdram_controller_0_s1_byteenable;                       // mm_interconnect_1:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire         mm_interconnect_1_new_sdram_controller_0_s1_readdatavalid;                    // new_sdram_controller_0:za_valid -> mm_interconnect_1:new_sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_1_new_sdram_controller_0_s1_write;                            // mm_interconnect_1:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire  [15:0] mm_interconnect_1_new_sdram_controller_0_s1_writedata;                        // mm_interconnect_1:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire         mm_interconnect_1_audio_0_avalon_audio_slave_chipselect;                      // mm_interconnect_1:audio_0_avalon_audio_slave_chipselect -> audio_0:chipselect
	wire  [31:0] mm_interconnect_1_audio_0_avalon_audio_slave_readdata;                        // audio_0:readdata -> mm_interconnect_1:audio_0_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_1_audio_0_avalon_audio_slave_address;                         // mm_interconnect_1:audio_0_avalon_audio_slave_address -> audio_0:address
	wire         mm_interconnect_1_audio_0_avalon_audio_slave_read;                            // mm_interconnect_1:audio_0_avalon_audio_slave_read -> audio_0:read
	wire         mm_interconnect_1_audio_0_avalon_audio_slave_write;                           // mm_interconnect_1:audio_0_avalon_audio_slave_write -> audio_0:write
	wire  [31:0] mm_interconnect_1_audio_0_avalon_audio_slave_writedata;                       // mm_interconnect_1:audio_0_avalon_audio_slave_writedata -> audio_0:writedata
	wire  [31:0] mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_readdata;   // video_dma_controller_0:slave_readdata -> mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_address;    // mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_address -> video_dma_controller_0:slave_address
	wire         mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_read;       // mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_read -> video_dma_controller_0:slave_read
	wire   [3:0] mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_byteenable; // mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_byteenable -> video_dma_controller_0:slave_byteenable
	wire         mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_write;      // mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_write -> video_dma_controller_0:slave_write
	wire  [31:0] mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_writedata;  // mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_writedata -> video_dma_controller_0:slave_writedata
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect;                   // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata;                     // jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest;                  // jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address;                      // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;                         // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;                        // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata;                    // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_1_nios2_qsys_0_debug_mem_slave_readdata;                      // nios2_qsys_0:debug_mem_slave_readdata -> mm_interconnect_1:nios2_qsys_0_debug_mem_slave_readdata
	wire         mm_interconnect_1_nios2_qsys_0_debug_mem_slave_waitrequest;                   // nios2_qsys_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_qsys_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_1_nios2_qsys_0_debug_mem_slave_debugaccess;                   // mm_interconnect_1:nios2_qsys_0_debug_mem_slave_debugaccess -> nios2_qsys_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_1_nios2_qsys_0_debug_mem_slave_address;                       // mm_interconnect_1:nios2_qsys_0_debug_mem_slave_address -> nios2_qsys_0:debug_mem_slave_address
	wire         mm_interconnect_1_nios2_qsys_0_debug_mem_slave_read;                          // mm_interconnect_1:nios2_qsys_0_debug_mem_slave_read -> nios2_qsys_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_1_nios2_qsys_0_debug_mem_slave_byteenable;                    // mm_interconnect_1:nios2_qsys_0_debug_mem_slave_byteenable -> nios2_qsys_0:debug_mem_slave_byteenable
	wire         mm_interconnect_1_nios2_qsys_0_debug_mem_slave_write;                         // mm_interconnect_1:nios2_qsys_0_debug_mem_slave_write -> nios2_qsys_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_1_nios2_qsys_0_debug_mem_slave_writedata;                     // mm_interconnect_1:nios2_qsys_0_debug_mem_slave_writedata -> nios2_qsys_0:debug_mem_slave_writedata
	wire         mm_interconnect_1_onchip_memory2_0_s1_chipselect;                             // mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_readdata;                               // onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	wire  [10:0] mm_interconnect_1_onchip_memory2_0_s1_address;                                // mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_1_onchip_memory2_0_s1_byteenable;                             // mm_interconnect_1:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_1_onchip_memory2_0_s1_write;                                  // mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_writedata;                              // mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_1_onchip_memory2_0_s1_clken;                                  // mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver0_irq;                                                     // audio_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                     // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_qsys_0_irq_irq;                                                         // irq_mapper:sender_irq -> nios2_qsys_0:irq
	wire         rst_controller_reset_out_reset;                                               // rst_controller:reset_out -> [audio_0:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_1:nios2_qsys_0_reset_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, nios2_qsys_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                           // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                           // rst_controller_001:reset_out -> [mm_interconnect_0:avalon_MM_4_to_1_adapter_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:video_dma_controller_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:avalon_MM_4_to_1_adapter_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:video_dma_controller_0_reset_reset_bridge_in_reset_reset, video_dma_controller_0:reset, video_vga_controller_0:reset]

	sub_top_audio_0 audio_0 (
		.clk         (sys_sdram_pll_0_sdram_clk_clk),                           //                clk.clk
		.reset       (rst_controller_reset_out_reset),                          //              reset.reset
		.address     (mm_interconnect_1_audio_0_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_1_audio_0_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_1_audio_0_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_1_audio_0_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_1_audio_0_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_1_audio_0_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver0_irq),                                //          interrupt.irq
		.AUD_BCLK    (audio_0_external_interface_BCLK),                         // external_interface.export
		.AUD_DACDAT  (audio_0_external_interface_DACDAT),                       //                   .export
		.AUD_DACLRCK (audio_0_external_interface_DACLRCK)                       //                   .export
	);

	avalon_MM_4_to_1_adapter avalon_mm_4_to_1_adapter_0 (
		.clock           (sys_sdram_pll_0_sys_clk_clk),                                             //   clock_reset.clk
		.reset_n         (~sys_sdram_pll_0_reset_source_reset),                                     //         reset.reset_n
		.m_waitrequest   (avalon_mm_4_to_1_adapter_0_avalon_master_waitrequest),                    // avalon_master.waitrequest
		.m_address       (avalon_mm_4_to_1_adapter_0_avalon_master_address),                        //              .address
		.m_byteenable    (avalon_mm_4_to_1_adapter_0_avalon_master_byteenable),                     //              .byteenable
		.m_read          (avalon_mm_4_to_1_adapter_0_avalon_master_read),                           //              .read
		.m_readdata      (avalon_mm_4_to_1_adapter_0_avalon_master_readdata),                       //              .readdata
		.m_readdatavalid (avalon_mm_4_to_1_adapter_0_avalon_master_readdatavalid),                  //              .readdatavalid
		.m_chipselect    (avalon_mm_4_to_1_adapter_0_avalon_master_chipselect),                     //              .chipselect
		.m_lock          (avalon_mm_4_to_1_adapter_0_avalon_master_lock),                           //              .lock
		.s_waitrequest   (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_waitrequest),   //  avalon_slave.waitrequest
		.s_readdata      (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_readdata),      //              .readdata
		.s_address       (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_address),       //              .address
		.s_read          (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_read),          //              .read
		.s_readdatavalid (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_readdatavalid), //              .readdatavalid
		.s_lock          (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_lock)           //              .lock
	);

	sub_top_jtag_uart_0 jtag_uart_0 (
		.clk            (sys_sdram_pll_0_sdram_clk_clk),                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	sub_top_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (sys_sdram_pll_0_sdram_clk_clk),                             //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                           // reset.reset_n
		.az_addr        (mm_interconnect_1_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (new_sdram_controller_0_wire_addr),                          //  wire.export
		.zs_ba          (new_sdram_controller_0_wire_ba),                            //      .export
		.zs_cas_n       (new_sdram_controller_0_wire_cas_n),                         //      .export
		.zs_cke         (new_sdram_controller_0_wire_cke),                           //      .export
		.zs_cs_n        (new_sdram_controller_0_wire_cs_n),                          //      .export
		.zs_dq          (new_sdram_controller_0_wire_dq),                            //      .export
		.zs_dqm         (new_sdram_controller_0_wire_dqm),                           //      .export
		.zs_ras_n       (new_sdram_controller_0_wire_ras_n),                         //      .export
		.zs_we_n        (new_sdram_controller_0_wire_we_n)                           //      .export
	);

	sub_top_nios2_qsys_0 nios2_qsys_0 (
		.clk                                 (sys_sdram_pll_0_sdram_clk_clk),                              //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_qsys_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_qsys_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	sub_top_onchip_memory2_0 onchip_memory2_0 (
		.clk        (sys_sdram_pll_0_sdram_clk_clk),                    //   clk1.clk
		.address    (mm_interconnect_1_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	sub_top_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n),                     //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sys_sdram_pll_0_sdram_clk_clk),      //    sdram_clk.clk
		.reset_source_reset (sys_sdram_pll_0_reset_source_reset)  // reset_source.reset
	);

	sub_top_video_dma_controller_0 video_dma_controller_0 (
		.clk                  (sys_sdram_pll_0_sys_clk_clk),                                                  //                      clk.clk
		.reset                (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.master_address       (video_dma_controller_0_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (video_dma_controller_0_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_arbiterlock   (video_dma_controller_0_avalon_dma_master_lock),                                //                         .lock
		.master_read          (video_dma_controller_0_avalon_dma_master_read),                                //                         .read
		.master_readdata      (video_dma_controller_0_avalon_dma_master_readdata),                            //                         .readdata
		.master_readdatavalid (video_dma_controller_0_avalon_dma_master_readdatavalid),                       //                         .readdatavalid
		.slave_address        (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_readdata),   //                         .readdata
		.stream_ready         (video_dma_controller_0_avalon_pixel_source_ready),                             //      avalon_pixel_source.ready
		.stream_data          (video_dma_controller_0_avalon_pixel_source_data),                              //                         .data
		.stream_startofpacket (video_dma_controller_0_avalon_pixel_source_startofpacket),                     //                         .startofpacket
		.stream_endofpacket   (video_dma_controller_0_avalon_pixel_source_endofpacket),                       //                         .endofpacket
		.stream_valid         (video_dma_controller_0_avalon_pixel_source_valid)                              //                         .valid
	);

	sub_top_video_vga_controller_0 video_vga_controller_0 (
		.clk           (sys_sdram_pll_0_sys_clk_clk),                              //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),                       //              reset.reset
		.data          (video_dma_controller_0_avalon_pixel_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dma_controller_0_avalon_pixel_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dma_controller_0_avalon_pixel_source_endofpacket),   //                   .endofpacket
		.valid         (video_dma_controller_0_avalon_pixel_source_valid),         //                   .valid
		.ready         (video_dma_controller_0_avalon_pixel_source_ready),         //                   .ready
		.VGA_CLK       (video_vga_controller_0_external_interface_CLK),            // external_interface.export
		.VGA_HS        (video_vga_controller_0_external_interface_HS),             //                   .export
		.VGA_VS        (video_vga_controller_0_external_interface_VS),             //                   .export
		.VGA_BLANK     (video_vga_controller_0_external_interface_BLANK),          //                   .export
		.VGA_SYNC      (video_vga_controller_0_external_interface_SYNC),           //                   .export
		.VGA_R         (video_vga_controller_0_external_interface_R),              //                   .export
		.VGA_G         (video_vga_controller_0_external_interface_G),              //                   .export
		.VGA_B         (video_vga_controller_0_external_interface_B)               //                   .export
	);

	sub_top_mm_interconnect_0 mm_interconnect_0 (
		.sys_sdram_pll_0_sys_clk_clk                                  (sys_sdram_pll_0_sys_clk_clk),                                             //                                sys_sdram_pll_0_sys_clk.clk
		.avalon_MM_4_to_1_adapter_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                      // avalon_MM_4_to_1_adapter_0_reset_reset_bridge_in_reset.reset
		.video_dma_controller_0_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                                      //     video_dma_controller_0_reset_reset_bridge_in_reset.reset
		.video_dma_controller_0_avalon_dma_master_address             (video_dma_controller_0_avalon_dma_master_address),                        //               video_dma_controller_0_avalon_dma_master.address
		.video_dma_controller_0_avalon_dma_master_waitrequest         (video_dma_controller_0_avalon_dma_master_waitrequest),                    //                                                       .waitrequest
		.video_dma_controller_0_avalon_dma_master_read                (video_dma_controller_0_avalon_dma_master_read),                           //                                                       .read
		.video_dma_controller_0_avalon_dma_master_readdata            (video_dma_controller_0_avalon_dma_master_readdata),                       //                                                       .readdata
		.video_dma_controller_0_avalon_dma_master_readdatavalid       (video_dma_controller_0_avalon_dma_master_readdatavalid),                  //                                                       .readdatavalid
		.video_dma_controller_0_avalon_dma_master_lock                (video_dma_controller_0_avalon_dma_master_lock),                           //                                                       .lock
		.avalon_MM_4_to_1_adapter_0_avalon_slave_address              (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_address),       //                avalon_MM_4_to_1_adapter_0_avalon_slave.address
		.avalon_MM_4_to_1_adapter_0_avalon_slave_read                 (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_read),          //                                                       .read
		.avalon_MM_4_to_1_adapter_0_avalon_slave_readdata             (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_readdata),      //                                                       .readdata
		.avalon_MM_4_to_1_adapter_0_avalon_slave_readdatavalid        (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_readdatavalid), //                                                       .readdatavalid
		.avalon_MM_4_to_1_adapter_0_avalon_slave_waitrequest          (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_waitrequest),   //                                                       .waitrequest
		.avalon_MM_4_to_1_adapter_0_avalon_slave_lock                 (mm_interconnect_0_avalon_mm_4_to_1_adapter_0_avalon_slave_lock)           //                                                       .lock
	);

	sub_top_mm_interconnect_1 mm_interconnect_1 (
		.sys_sdram_pll_0_sdram_clk_clk                                (sys_sdram_pll_0_sdram_clk_clk),                                                //                              sys_sdram_pll_0_sdram_clk.clk
		.sys_sdram_pll_0_sys_clk_clk                                  (sys_sdram_pll_0_sys_clk_clk),                                                  //                                sys_sdram_pll_0_sys_clk.clk
		.avalon_MM_4_to_1_adapter_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                           // avalon_MM_4_to_1_adapter_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                                               //               nios2_qsys_0_reset_reset_bridge_in_reset.reset
		.video_dma_controller_0_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                                           //     video_dma_controller_0_reset_reset_bridge_in_reset.reset
		.avalon_MM_4_to_1_adapter_0_avalon_master_address             (avalon_mm_4_to_1_adapter_0_avalon_master_address),                             //               avalon_MM_4_to_1_adapter_0_avalon_master.address
		.avalon_MM_4_to_1_adapter_0_avalon_master_waitrequest         (avalon_mm_4_to_1_adapter_0_avalon_master_waitrequest),                         //                                                       .waitrequest
		.avalon_MM_4_to_1_adapter_0_avalon_master_byteenable          (avalon_mm_4_to_1_adapter_0_avalon_master_byteenable),                          //                                                       .byteenable
		.avalon_MM_4_to_1_adapter_0_avalon_master_chipselect          (avalon_mm_4_to_1_adapter_0_avalon_master_chipselect),                          //                                                       .chipselect
		.avalon_MM_4_to_1_adapter_0_avalon_master_read                (avalon_mm_4_to_1_adapter_0_avalon_master_read),                                //                                                       .read
		.avalon_MM_4_to_1_adapter_0_avalon_master_readdata            (avalon_mm_4_to_1_adapter_0_avalon_master_readdata),                            //                                                       .readdata
		.avalon_MM_4_to_1_adapter_0_avalon_master_readdatavalid       (avalon_mm_4_to_1_adapter_0_avalon_master_readdatavalid),                       //                                                       .readdatavalid
		.avalon_MM_4_to_1_adapter_0_avalon_master_lock                (avalon_mm_4_to_1_adapter_0_avalon_master_lock),                                //                                                       .lock
		.nios2_qsys_0_data_master_address                             (nios2_qsys_0_data_master_address),                                             //                               nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                                         //                                                       .waitrequest
		.nios2_qsys_0_data_master_byteenable                          (nios2_qsys_0_data_master_byteenable),                                          //                                                       .byteenable
		.nios2_qsys_0_data_master_read                                (nios2_qsys_0_data_master_read),                                                //                                                       .read
		.nios2_qsys_0_data_master_readdata                            (nios2_qsys_0_data_master_readdata),                                            //                                                       .readdata
		.nios2_qsys_0_data_master_write                               (nios2_qsys_0_data_master_write),                                               //                                                       .write
		.nios2_qsys_0_data_master_writedata                           (nios2_qsys_0_data_master_writedata),                                           //                                                       .writedata
		.nios2_qsys_0_data_master_debugaccess                         (nios2_qsys_0_data_master_debugaccess),                                         //                                                       .debugaccess
		.nios2_qsys_0_instruction_master_address                      (nios2_qsys_0_instruction_master_address),                                      //                        nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest                  (nios2_qsys_0_instruction_master_waitrequest),                                  //                                                       .waitrequest
		.nios2_qsys_0_instruction_master_read                         (nios2_qsys_0_instruction_master_read),                                         //                                                       .read
		.nios2_qsys_0_instruction_master_readdata                     (nios2_qsys_0_instruction_master_readdata),                                     //                                                       .readdata
		.audio_0_avalon_audio_slave_address                           (mm_interconnect_1_audio_0_avalon_audio_slave_address),                         //                             audio_0_avalon_audio_slave.address
		.audio_0_avalon_audio_slave_write                             (mm_interconnect_1_audio_0_avalon_audio_slave_write),                           //                                                       .write
		.audio_0_avalon_audio_slave_read                              (mm_interconnect_1_audio_0_avalon_audio_slave_read),                            //                                                       .read
		.audio_0_avalon_audio_slave_readdata                          (mm_interconnect_1_audio_0_avalon_audio_slave_readdata),                        //                                                       .readdata
		.audio_0_avalon_audio_slave_writedata                         (mm_interconnect_1_audio_0_avalon_audio_slave_writedata),                       //                                                       .writedata
		.audio_0_avalon_audio_slave_chipselect                        (mm_interconnect_1_audio_0_avalon_audio_slave_chipselect),                      //                                                       .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                        (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),                      //                          jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                          (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),                        //                                                       .write
		.jtag_uart_0_avalon_jtag_slave_read                           (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),                         //                                                       .read
		.jtag_uart_0_avalon_jtag_slave_readdata                       (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),                     //                                                       .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                      (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),                    //                                                       .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                    (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest),                  //                                                       .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),                   //                                                       .chipselect
		.new_sdram_controller_0_s1_address                            (mm_interconnect_1_new_sdram_controller_0_s1_address),                          //                              new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                              (mm_interconnect_1_new_sdram_controller_0_s1_write),                            //                                                       .write
		.new_sdram_controller_0_s1_read                               (mm_interconnect_1_new_sdram_controller_0_s1_read),                             //                                                       .read
		.new_sdram_controller_0_s1_readdata                           (mm_interconnect_1_new_sdram_controller_0_s1_readdata),                         //                                                       .readdata
		.new_sdram_controller_0_s1_writedata                          (mm_interconnect_1_new_sdram_controller_0_s1_writedata),                        //                                                       .writedata
		.new_sdram_controller_0_s1_byteenable                         (mm_interconnect_1_new_sdram_controller_0_s1_byteenable),                       //                                                       .byteenable
		.new_sdram_controller_0_s1_readdatavalid                      (mm_interconnect_1_new_sdram_controller_0_s1_readdatavalid),                    //                                                       .readdatavalid
		.new_sdram_controller_0_s1_waitrequest                        (mm_interconnect_1_new_sdram_controller_0_s1_waitrequest),                      //                                                       .waitrequest
		.new_sdram_controller_0_s1_chipselect                         (mm_interconnect_1_new_sdram_controller_0_s1_chipselect),                       //                                                       .chipselect
		.nios2_qsys_0_debug_mem_slave_address                         (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_address),                       //                           nios2_qsys_0_debug_mem_slave.address
		.nios2_qsys_0_debug_mem_slave_write                           (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_write),                         //                                                       .write
		.nios2_qsys_0_debug_mem_slave_read                            (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_read),                          //                                                       .read
		.nios2_qsys_0_debug_mem_slave_readdata                        (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_readdata),                      //                                                       .readdata
		.nios2_qsys_0_debug_mem_slave_writedata                       (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_writedata),                     //                                                       .writedata
		.nios2_qsys_0_debug_mem_slave_byteenable                      (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_byteenable),                    //                                                       .byteenable
		.nios2_qsys_0_debug_mem_slave_waitrequest                     (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_waitrequest),                   //                                                       .waitrequest
		.nios2_qsys_0_debug_mem_slave_debugaccess                     (mm_interconnect_1_nios2_qsys_0_debug_mem_slave_debugaccess),                   //                                                       .debugaccess
		.onchip_memory2_0_s1_address                                  (mm_interconnect_1_onchip_memory2_0_s1_address),                                //                                    onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                    (mm_interconnect_1_onchip_memory2_0_s1_write),                                  //                                                       .write
		.onchip_memory2_0_s1_readdata                                 (mm_interconnect_1_onchip_memory2_0_s1_readdata),                               //                                                       .readdata
		.onchip_memory2_0_s1_writedata                                (mm_interconnect_1_onchip_memory2_0_s1_writedata),                              //                                                       .writedata
		.onchip_memory2_0_s1_byteenable                               (mm_interconnect_1_onchip_memory2_0_s1_byteenable),                             //                                                       .byteenable
		.onchip_memory2_0_s1_chipselect                               (mm_interconnect_1_onchip_memory2_0_s1_chipselect),                             //                                                       .chipselect
		.onchip_memory2_0_s1_clken                                    (mm_interconnect_1_onchip_memory2_0_s1_clken),                                  //                                                       .clken
		.video_dma_controller_0_avalon_dma_control_slave_address      (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_address),    //        video_dma_controller_0_avalon_dma_control_slave.address
		.video_dma_controller_0_avalon_dma_control_slave_write        (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_write),      //                                                       .write
		.video_dma_controller_0_avalon_dma_control_slave_read         (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_read),       //                                                       .read
		.video_dma_controller_0_avalon_dma_control_slave_readdata     (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_readdata),   //                                                       .readdata
		.video_dma_controller_0_avalon_dma_control_slave_writedata    (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_writedata),  //                                                       .writedata
		.video_dma_controller_0_avalon_dma_control_slave_byteenable   (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_byteenable)  //                                                       .byteenable
	);

	sub_top_irq_mapper irq_mapper (
		.clk           (sys_sdram_pll_0_sdram_clk_clk),  //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_qsys_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (sys_sdram_pll_0_reset_source_reset), // reset_in0.reset
		.clk            (sys_sdram_pll_0_sdram_clk_clk),      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (sys_sdram_pll_0_reset_source_reset), // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
